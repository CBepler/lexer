module simple_logic (
    input wire a,
    output wire b, //Comment
);
endmodule
